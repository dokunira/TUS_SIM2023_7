*SUBCKT Definition - CMOS INVERTER -

* 1:in 2:out 3:Vdd
.SUBCKT Schmitt_INV 1 2 3

*M Drain Gate Source BackSource ModelName
MP1 4 1 3 3 pmos1
MP2 2 1 4 3 pmos1
MP3 0 2 4 3 pmos1
MN1 2 1 5 0 nmos1
MN2 5 1 0 0 nmos1 
MN3 3 2 0 0 nmos1

*parasitic capacitance
CL 2 0 0.05p

.ENDS