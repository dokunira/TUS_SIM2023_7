TEST DFF

.INCLUDE DFF.cir

*.MODEL モデル名 タイプ(パラメータ1 = パラメータ値1 …)
*level:モデル番号 vto:閾値電圧 l:チャネル長 w:チャネル幅 tox:酸化膜の厚さ cbd:BD間寄生容量 cbs:BS間寄生容量
* .MODEL nmos1 nmos(level=3 vto=1 l=1u w=10u tox=0.5u cbd=20f cbs=20f)
* .MODEL pmos1 pmos(level=3 vto=-1 l=1u w=10u tox=0.5u cbd=20f cbs=20f)
.MODEL nmos1 nmos(vto=1)
.MODEL pmos1 pmos(vto=-1)

* 1:D 2:CK 3:Q 4:invQ 5:Vdd DFF
X1 1 2 3 4 5 DFF

VCC 5 0 DC=5
* PWL(時間 値 時間 値 ・・・)
VD 1 0 PWL(0 0 0.9u 0 1u 5 3u 5 3.1u 0 6u 0 6.1u 5 10u 5)
* PULSE(初期値 波高値 遅延時間 立上がり時間 立下り時間 パルス幅 周期)
VCK 2 0 PULSE(0 5 0.5u 50n 50n 1u 2u)

*.TRAN 刻み 終了時刻
.TRAN 1n 10u
.END